module module_s(input logic a,b, output logic y1);

and U1 (y1,a,b);

// Complete for OR and XOR gates

endmodule
